`define REG_R0 4'h0
`define REG_R1 4'h1
`define REG_R2 4'h2
`define REG_R3 4'h3
`define REG_R4 4'h4
`define REG_R5 4'h5
`define REG_R6 4'h6
`define REG_R7 4'h7
`define REG_R8 4'h8
`define REG_R9 4'h9
`define REG_R10 4'ha
`define REG_R11 4'hb
`define REG_R12 4'hc
`define REG_PC 4'hd
`define REG_SP 4'he
`define REG_FP 4'hf
