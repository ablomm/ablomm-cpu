module cu_tb;
  import cpu_pkg::*;
  import reg_pkg::*;

  logic clk;
  logic start;
  logic hwint;
  logic rst = 0;
  ir_t ir_value;
  status_t status_value;

  // control signals
  logic mem_rd;
  logic mem_wr;

  logic oe_alu;
  logic [3:0] alu_op;

  logic [31:0] a_reg_mask;
  logic [31:0] b_reg_mask;

  reg_e sel_a_reg;
  reg_e sel_b_reg;
  reg_e sel_in_reg;

  logic oe_a_reg_file;
  logic oe_b_reg_file;
  logic ld_reg_file;
  logic post_inc_sp;
  logic pre_dec_sp;
  logic post_inc_pc;

  logic oe_a_consts;
  logic oe_b_consts;

  logic oe_a_ir;
  logic oe_b_ir;
  logic ld_ir;

  logic ld_alu_status;
  logic imask_in;
  logic ld_imask;
  cpu_mode_e mode_in;
  logic ld_mode;

  cu cu0 (
      .*,
      .ir(ir_value),
      .status(status_value)
  );


  initial begin
    // STOP state
    clk = 0;
    #1;

    start = 1;
    clk   = 1;
    #1;

    // FETCH state
    clk = 0;
    #1;
    $display("sel_b_reg: %d, oe_b_reg_file: %d, mem_rd: %d, ld_ir: %d, post_inc_pc: %d", sel_b_reg,
             oe_b_reg_file, mem_rd, ld_ir, post_inc_pc);

    assert (sel_b_reg === reg_pkg::PC && oe_b_reg_file === 1 && mem_rd === 1 && post_inc_pc === 1);
    clk = 1;
    start = 0;
    ir_value.condition = NONE;
    ir_value.instruction = alu_pkg::AND;
    ir_value.params.alu_op.flags.immediate = 0;
    ir_value.params.alu_op.flags.reverse = 0;
    ir_value.params.alu_op.flags.load = 1;
    ir_value.params.alu_op.flags.set_status = 0;
    ir_value.params.alu_op.reg_a = reg_pkg::R0;
    ir_value.params.alu_op.reg_b = reg_pkg::R1;
    ir_value.params.alu_op.reg_c = reg_pkg::R2;
    #1;

    // AND state
    clk = 0;
    #1;
    $display(
        "sel_a_reg: %d, oe_a_reg_file: %d, sel_b_reg: %d, oe_b_reg_file: %d, alu_op: %d, sel_in_reg: %d, ld_reg_file: %d",
        sel_a_reg, oe_a_reg_file, sel_b_reg, oe_b_reg_file, alu_op, sel_in_reg, ld_reg_file);

    assert (sel_a_reg === reg_pkg::R1 && oe_a_reg_file === 1 && sel_b_reg === reg_pkg::R2 && oe_b_reg_file === 1 && alu_op === alu_pkg::AND && sel_in_reg === reg_pkg::R0 && ld_reg_file === 1);
    clk = 1;
  end
endmodule
