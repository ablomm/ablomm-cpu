`define ALU_PASSA 4'h0
`define ALU_PASSB 4'h1

`define ALU_AND 4'h2
`define ALU_OR 4'h3
`define ALU_XOR 4'h4
`define ALU_NOT 4'h5

`define ALU_ADD 4'h6
`define ALU_ADDC 4'h7
`define ALU_SUB 4'h8
`define ALU_SUBB 4'h9
`define ALU_SHL 4'ha
`define ALU_SHR 4'hb
`define ALU_ASHR 4'hc
