import alu_pkg::*;
import reg_pkg::*;

module alu (
    input oe,
    input alu_op_e operation,
    input carry_in,
    input [31:0] a,
    input [31:0] b,
    output tri [31:0] out,
    output alu_status_t status
);

  logic [31:0] out_reg;

  assign out = oe ? out_reg : 'hz;

  always_comb begin
    case (operation)
      alu_pkg::PASSA: out_reg = a;
      alu_pkg::PASSB: out_reg = b;

      alu_pkg::AND: out_reg = a & b;
      alu_pkg::OR:  out_reg = a | b;
      alu_pkg::XOR: out_reg = a ^ b;
      alu_pkg::NOT: out_reg = ~a;

      alu_pkg::ADD: {status.carry, out_reg} = a + b;
      alu_pkg::ADDC: {status.carry, out_reg} = a + b + carry_in;
      alu_pkg::SUB: {status.carry, out_reg} = a - b;
      alu_pkg::SUBB: {status.carry, out_reg} = a - b - ~carry_in;
      alu_pkg::SHL: {status.carry, out_reg} = a << b;
      alu_pkg::SHR: out_reg = a >> b;
      alu_pkg::ASHR: out_reg = a >>> b;
      default: out_reg = 0;
    endcase
  end

  always @(out_reg) begin
    // negative
    status.negative = out_reg[31];

    // zero
    status.zero = out_reg === 0;

    // overflow
    status.overflow = out_reg[31] ^ a[31] ^ b[31] ^ status.carry;
  end
endmodule
